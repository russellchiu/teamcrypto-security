`ifndef CONSTANTS
`define CONSTANTS 1
// Constants
`define key_size 80
// `define key_size 128;
`define size 64
`define num_rounds 32

// sizes are defined for the blocks that are used
`define BLOCKSIZE 4
`define ARRSIZE 16
`endif

`define num_vectors 20
`define counter_bits 5

module Test_Constants();

endmodule
